`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:  Team Zigma
// Engineer: Nuwan Udara
// 
// Create Date: 31.01.2023 18:07:12
// Design Name: 
// Module Name: inDecode
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////



module inDecode(
    input 	   [31:0] inst,
    output reg [6:0] opcode,  
    output reg [4:0] rsAddr, //rs1
    output reg [4:0] rdAddr, //rd
    output reg [4:0] shamt,  //SHIFT VAL AND RS2
    output reg [3:0] alu_func,   // FOR ALU_contoller func_3 + 1 bit for add sub chnage like things
    output reg [31:0] imm,   // i TYPE  imm
    output reg [31:0] label // for braching
    );

always @(*)
	begin
	opcode=inst[31:25];       //Opcode is always the first 7 bits
	
	if(opcode==7'b0110011)        //Arithmetic and Shift Operations
		begin
		rsAddr<=  inst[16:12];
		rdAddr<=  inst[24:20];
		shamt<=   inst[11:7];
		alu_func<={inst[1],inst[19:17]}; //only for R instructions need inst[1],0
		imm<=32'b0;          
		label<=32'b0;
		end

	else if(opcode==7'b0010011)   //Immediate Operations
		begin
		rsAddr<=inst[16:12];
		rdAddr<=inst[24:20];
		shamt<=5'b00000;     // no need second address
		alu_func<={1'b0,inst[19:17]}; // no need for a sign bit from function 7
		imm<=inst[11:0];    
		label<=32'b0;   //only for U and UJ
		end
	else if(opcode==7'b0000011)   //Load Operations only using LW still pass function_3, this is basicly a I nstruction
		begin
		rsAddr<=inst[16:12]; //rs1
		rdAddr<=inst[24:20]; //rd
		shamt<=5'b00000;     // no need second address
		alu_func<={1'b0,inst[19:17]}; // no need for a sign bit from function 7
		imm<=inst[11:0];    //immediate value sign extended
		label<=32'b0;  	    // no need for this, only used in U and UJ
		end
    
    else if(opcode==7'b0100011)   //Store Operations Only Store Word, SW S instrucctions
		begin
		rsAddr<=inst[28:24];
		rdAddr<= 5'b00000;    //inst[23:19]; // will be used to take from the ALU result, if rdAddr =0, use write address from ALU result
		shamt<=5'b00000;      //no need this
		alu_func<={1'b0,inst[19:17]};
		imm<={inst[6:0],inst[24:20]};  // MSB and LSM in order
		label<=32'b0;   //No need this
		end

	else if(opcode==7'b1100011)    //Branch/Jump Operations   //BEQ, BLT, BLTU, BNE, SB; "B" instructions
		begin
		rsAddr<=inst[28:24]; // rs1 adddress
		rdAddr<=5'b0;
		shamt<=5'b0;
		alu_func<={1'b0,inst[19:17]};
		imm<={inst[0],inst[24],inst[6:1],inst[23:20],1'b0};   //{1'b0,inst[23:20],inst[6:1],inst[24],inst[0]}
		//label<=inst[28:4];
		label <= 32'b0;
		end

	else if(opcode==7'b1101111)    //J - JAL
		begin
		rsAddr<=5'b0;
		rdAddr<=5'b0;
		shamt<=5'b0;

		alu_func<=4'b0;
		imm<=32'b0;
		label<={inst[0],inst[19:12],imm[11],imm[10:1],1'b0}; // will be sign extended
		end

    else if(opcode==7'b1100111)    //I-type  JALR
		begin
		rsAddr<=inst[16:12];
		rdAddr<=inst[24:20];
		shamt<=5'b00000;     // no need second address
		alu_func<={1'b0,inst[19:17]}; // no need for a sign bit from function 7
		imm<=inst[11:0];
		label<=32'b0;
		end
    
    else if(opcode==7'b0110111)    //Upper LUI
		begin
		rsAddr<=5'b0;
		rdAddr<=inst[24:20];
		shamt<=5'b0;
		alu_func<=4'b0;
		imm<=32'b0;
		label<={inst[19:0],12'b0};
		end
    
    else if(opcode==7'b0010111)    //Upper AUIPC
		begin
		rsAddr<=5'b0;
		rdAddr<=inst[24:20];
		shamt<=5'b0;
		alu_func<=4'b0;
		imm<=32'b0;
		label<={inst[19:0],12'b0};
		end


	else                 //invalid instruction/empty instruction: make everything 0
		begin
		rsAddr<=5'b0;
		rdAddr<=5'b0;
		shamt<=5'b0;
		alu_func<=4'b0;
		imm<=32'b0;
		label<=32'b0;
		end
	end

// always @(*)                 //Assign MemWrite
// 	begin
// 		if(opcode==3'd2 & alu_func==4'd1)   //only in case of store word make it 1 ?
// 			begin
// 			MemWrite<=1;
// 			end
// 		else
// 			MemWrite<=0;
// 	end
endmodule